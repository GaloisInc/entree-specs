(* Top-level Coq module that re-exports everything for clients of the library *)

From EnTree Require Export
     Basics.HeterogeneousRelations
     Basics.QuantType
     Basics.PolyList
     Core.EnTreeDefinition
     Core.SubEvent
     Eq.Eqit
     Ref.Padded
     Ref.EnTreeSpecDefinition
     Ref.MRecSpec
     Ref.SpecM
     Ref.LetRecRefines
     Ref.DefRefines
.
